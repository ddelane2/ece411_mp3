library verilog;
use verilog.vl_types.all;
entity nzpcomp_sv_unit is
end nzpcomp_sv_unit;
