library verilog;
use verilog.vl_types.all;
entity rom_control_sv_unit is
end rom_control_sv_unit;
