library verilog;
use verilog.vl_types.all;
entity if_id_ff_sv_unit is
end if_id_ff_sv_unit;
