library verilog;
use verilog.vl_types.all;
entity adju_sv_unit is
end adju_sv_unit;
