library verilog;
use verilog.vl_types.all;
entity id_ex_ff_sv_unit is
end id_ex_ff_sv_unit;
